	// Verilator lint_off UNUSED
	// These defined primitives are BIG_ENDIAN.  The first byte out is on
	// the left.  The first bit out is the LSB on the right.

				// Byte 0,	Byte 1,		Byte 2,		Byte 3
				// K.3b.5b,	D.3b.5b,	D.3b.5b,	D.3b.5b
				// Z.HGF.EDCBA
	localparam	[32:0]	P_ALIGN  = { 1'b1, 8'b101_11100, 8'b010_01010, 8'b010_01010, 8'b011_11011 },	// bc4a4a7b
				P_CONT   = { 1'b1, 8'b011_11100, 8'b101_01010, 8'b100_11001, 8'b100_11001 },	// 7caa9999
				P_DMAT   = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b001_10110, 8'b001_10110 },	// 7cb53636
				P_EOF    = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b110_10101, 8'b110_10101 },	// 7cb5d5d5
				P_HOLD   = { 1'b1, 8'b011_11100, 8'b101_01010, 8'b110_10101, 8'b110_10101 },	// 7caad5d5
				P_HOLDA  = { 1'b1, 8'b011_11100, 8'b101_01010, 8'b100_10101, 8'b100_10101 },	// 7caa9595
				P_PMACK  = { 1'b1, 8'b011_11100, 8'b100_10101, 8'b100_10101, 8'b100_10101 },	// 7c959595
				P_PMNAK  = { 1'b1, 8'b011_11100, 8'b100_10101, 8'b111_10101, 8'b111_10101 },	// 7c95f5f5
				P_PMREQ_P= { 1'b1, 8'b011_11100, 8'b101_10101, 8'b000_10111, 8'b000_10111 },	// 7cb51717
				P_PMREQ_S= { 1'b1, 8'b011_11100, 8'b100_10101, 8'b011_10101, 8'b011_10101 },	// 7c957575
				P_R_ERR  = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b010_10110, 8'b010_10110 },	// 7cb55656
				P_R_IP   = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b010_10101, 8'b010_10101 },	// 7cb55555
				P_R_OK   = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b001_10101, 8'b001_10101 },	// 7cb53535
				P_R_RDY  = { 1'b1, 8'b011_11100, 8'b100_10101, 8'b010_01010, 8'b010_01010 },	// 7c954a4a
				P_SOF    = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b001_10111, 8'b001_10111 },	// 7cb53737
				P_SYNC   = { 1'b1, 8'b011_11100, 8'b100_10101, 8'b101_10101, 8'b101_10101 },	// 7c95b5b5
				P_WTRM   = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b010_11000, 8'b010_11000 },	// 7cb55858
				P_X_RDY  = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b010_10111, 8'b010_10111 },	// 7cb55757
				D10_2	 = 33'h04A4A4A4A;
	// Verilator lint_on  UNUSED
