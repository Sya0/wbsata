////////////////////////////////////////////////////////////////////////////////
//
// Filename:	bench/verilog/mdl_s10b8b.v
// {{{
// Project:	A Wishbone SATA controller
//
// Purpose:	An 8B/10B Decoder: receives 10bits at a time, produces 8bits
//		at the output.  Protocols are only nominally AXI Stream based.
//
// Creator:	Dan Gisselquist, Ph.D.
//		Gisselquist Technology, LLC
//
////////////////////////////////////////////////////////////////////////////////
// }}}
// Copyright (C) 2022-2025, Gisselquist Technology, LLC
// {{{
// This file is part of the WBSATA project.
//
// The WBSATA project is a free software (firmware) project: you may
// redistribute it and/or modify it under the terms of  the GNU General Public
// License as published by the Free Software Foundation, either version 3 of
// the License, or (at your option) any later version.
//
// This program is distributed in the hope that it will be useful, but WITHOUT
// ANY WARRANTY; without even the implied warranty of MERCHANTIBILITY or
// FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
// for more details.
//
// You should have received a copy of the GNU General Public License along
// with this program.  If not, please see <http://www.gnu.org/licenses/> for a
// copy.
// }}}
// License:	GPL, v3, as defined and found on www.gnu.org,
// {{{
//		http://www.gnu.org/licenses/gpl.html
//
////////////////////////////////////////////////////////////////////////////////
//
`default_nettype none
`timescale	1ns/1ps
// }}}
module	mdl_s10b8b (
		input	wire	[9:0]	S_DATA,
		//
		output	wire	[8:0]	M_DATA
	);

	//
	// decoded = XTRA, 5D, 3D
	//
	reg	[8:0]	decoded;
	wire	[5:0]	abcdei = S_DATA[9:4];
	wire	[3:0]	fghj   = S_DATA[3:0];

	always @(*)
	case({ abcdei, fghj })
	{ 6'b100_111, 4'b0100 }: decoded = { 1'b0, 5'd00, 3'h0 };	// RD-
	{ 6'b011_000, 4'b1011 }: decoded = { 1'b0, 5'd00, 3'h0 };	// RD+
	{ 6'b011_101, 4'b0100 }: decoded = { 1'b0, 5'd01, 3'h0 };	// RD-
	{ 6'b100_010, 4'b1011 }: decoded = { 1'b0, 5'd01, 3'h0 };	// RD+
	{ 6'b101_101, 4'b0100 }: decoded = { 1'b0, 5'd02, 3'h0 };	// RD-
	{ 6'b010_010, 4'b1011 }: decoded = { 1'b0, 5'd02, 3'h0 };	// RD+
	{ 6'b110_001, 4'b1011 }: decoded = { 1'b0, 5'd03, 3'h0 };	// RD-
	{ 6'b110_001, 4'b0100 }: decoded = { 1'b0, 5'd03, 3'h0 };	// RD+
	{ 6'b110_101, 4'b0100 }: decoded = { 1'b0, 5'd04, 3'h0 };	// RD-
	{ 6'b001_010, 4'b1011 }: decoded = { 1'b0, 5'd04, 3'h0 };	// RD+
	{ 6'b101_001, 4'b1011 }: decoded = { 1'b0, 5'd05, 3'h0 };	// RD-
	{ 6'b101_001, 4'b0100 }: decoded = { 1'b0, 5'd05, 3'h0 };	// RD+
	{ 6'b011_001, 4'b1011 }: decoded = { 1'b0, 5'd06, 3'h0 };	// RD-
	{ 6'b011_001, 4'b0100 }: decoded = { 1'b0, 5'd06, 3'h0 };	// RD+
	{ 6'b111_000, 4'b1011 }: decoded = { 1'b0, 5'd07, 3'h0 };	// RD-
	{ 6'b000_111, 4'b0100 }: decoded = { 1'b0, 5'd07, 3'h0 };	// RD+
	//
	{ 6'b111_001, 4'b0100 }: decoded = { 1'b0, 5'd08, 3'h0 };	// RD-
	{ 6'b000_110, 4'b1011 }: decoded = { 1'b0, 5'd08, 3'h0 };	// RD+
	{ 6'b100_101, 4'b1011 }: decoded = { 1'b0, 5'd09, 3'h0 };	// RD-
	{ 6'b100_101, 4'b0100 }: decoded = { 1'b0, 5'd09, 3'h0 };	// RD+
	{ 6'b010_101, 4'b1011 }: decoded = { 1'b0, 5'd10, 3'h0 };	// RD-
	{ 6'b010_101, 4'b0100 }: decoded = { 1'b0, 5'd10, 3'h0 };	// RD+
	{ 6'b110_100, 4'b1011 }: decoded = { 1'b0, 5'd11, 3'h0 };	// RD-
	{ 6'b110_100, 4'b0100 }: decoded = { 1'b0, 5'd11, 3'h0 };	// RD+
	{ 6'b001_101, 4'b1011 }: decoded = { 1'b0, 5'd12, 3'h0 };	// RD-
	{ 6'b001_101, 4'b0100 }: decoded = { 1'b0, 5'd12, 3'h0 };	// RD+
	{ 6'b101_100, 4'b1011 }: decoded = { 1'b0, 5'd13, 3'h0 };	// RD-
	{ 6'b101_100, 4'b0100 }: decoded = { 1'b0, 5'd13, 3'h0 };	// RD+
	{ 6'b011_100, 4'b1011 }: decoded = { 1'b0, 5'd14, 3'h0 };	// RD-
	{ 6'b011_100, 4'b0100 }: decoded = { 1'b0, 5'd14, 3'h0 };	// RD+
	{ 6'b010_111, 4'b0100 }: decoded = { 1'b0, 5'd15, 3'h0 };	// RD-
	{ 6'b101_000, 4'b1011 }: decoded = { 1'b0, 5'd15, 3'h0 };	// RD+
	//
	{ 6'b011_011, 4'b0100 }: decoded = { 1'b0, 5'd16, 3'h0 };	// RD-
	{ 6'b100_100, 4'b1011 }: decoded = { 1'b0, 5'd16, 3'h0 };	// RD+
	{ 6'b100_011, 4'b1011 }: decoded = { 1'b0, 5'd17, 3'h0 };	// RD-
	{ 6'b100_011, 4'b0100 }: decoded = { 1'b0, 5'd17, 3'h0 };	// RD+
	{ 6'b010_011, 4'b1011 }: decoded = { 1'b0, 5'd18, 3'h0 };	// RD-
	{ 6'b010_011, 4'b0100 }: decoded = { 1'b0, 5'd18, 3'h0 };	// RD+
	{ 6'b110_010, 4'b1011 }: decoded = { 1'b0, 5'd19, 3'h0 };	// RD-
	{ 6'b110_010, 4'b0100 }: decoded = { 1'b0, 5'd19, 3'h0 };	// RD+
	{ 6'b001_011, 4'b1011 }: decoded = { 1'b0, 5'd20, 3'h0 };	// RD-
	{ 6'b001_011, 4'b0100 }: decoded = { 1'b0, 5'd20, 3'h0 };	// RD+
	{ 6'b101_010, 4'b1011 }: decoded = { 1'b0, 5'd21, 3'h0 };	// RD-
	{ 6'b101_010, 4'b0100 }: decoded = { 1'b0, 5'd21, 3'h0 };	// RD+
	{ 6'b011_010, 4'b1011 }: decoded = { 1'b0, 5'd22, 3'h0 };	// RD-
	{ 6'b011_010, 4'b0100 }: decoded = { 1'b0, 5'd22, 3'h0 };	// RD+
	{ 6'b111_010, 4'b0100 }: decoded = { 1'b0, 5'd23, 3'h0 };	// RD-
	{ 6'b000_101, 4'b1011 }: decoded = { 1'b0, 5'd23, 3'h0 };	// RD+
	//
	{ 6'b110_011, 4'b0100 }: decoded = { 1'b0, 5'd24, 3'h0 };	// RD-
	{ 6'b001_100, 4'b1011 }: decoded = { 1'b0, 5'd24, 3'h0 };	// RD+
	{ 6'b100_110, 4'b1011 }: decoded = { 1'b0, 5'd25, 3'h0 };	// RD-
	{ 6'b100_110, 4'b0100 }: decoded = { 1'b0, 5'd25, 3'h0 };	// RD+
	{ 6'b010_110, 4'b1011 }: decoded = { 1'b0, 5'd26, 3'h0 };	// RD-
	{ 6'b010_110, 4'b0100 }: decoded = { 1'b0, 5'd26, 3'h0 };	// RD+
	{ 6'b110_110, 4'b0100 }: decoded = { 1'b0, 5'd27, 3'h0 };	// RD-
	{ 6'b001_001, 4'b1011 }: decoded = { 1'b0, 5'd27, 3'h0 };	// RD+
	{ 6'b001_110, 4'b1011 }: decoded = { 1'b0, 5'd28, 3'h0 };	// RD-
	{ 6'b001_110, 4'b0100 }: decoded = { 1'b0, 5'd28, 3'h0 };	// RD+
	{ 6'b101_110, 4'b0100 }: decoded = { 1'b0, 5'd29, 3'h0 };	// RD-
	{ 6'b010_001, 4'b1011 }: decoded = { 1'b0, 5'd29, 3'h0 };	// RD+
	{ 6'b011_110, 4'b0100 }: decoded = { 1'b0, 5'd30, 3'h0 };	// RD-
	{ 6'b100_001, 4'b1011 }: decoded = { 1'b0, 5'd30, 3'h0 };	// RD+
	{ 6'b101_011, 4'b0100 }: decoded = { 1'b0, 5'd31, 3'h0 };	// RD-
	{ 6'b010_100, 4'b1011 }: decoded = { 1'b0, 5'd31, 3'h0 };	// RD+
	//
	//
	//
	{ 6'b100_111, 4'b1001 }: decoded = { 1'b0, 5'd00, 3'h1 };	// RD-
	{ 6'b011_000, 4'b1001 }: decoded = { 1'b0, 5'd00, 3'h1 };	// RD+
	{ 6'b011_101, 4'b1001 }: decoded = { 1'b0, 5'd01, 3'h1 };	// RD-
	{ 6'b100_010, 4'b1001 }: decoded = { 1'b0, 5'd01, 3'h1 };	// RD+
	{ 6'b101_101, 4'b1001 }: decoded = { 1'b0, 5'd02, 3'h1 };	// RD-
	{ 6'b010_010, 4'b1001 }: decoded = { 1'b0, 5'd02, 3'h1 };	// RD+
	{ 6'b110_001, 4'b1001 }: decoded = { 1'b0, 5'd03, 3'h1 };	// RD-/+
	// { 6'b110_001, 4'b1001 }: decoded = { 1'b0, 5'd03, 3'h1 };	// RD+
	{ 6'b110_101, 4'b1001 }: decoded = { 1'b0, 5'd04, 3'h1 };	// RD-
	{ 6'b001_010, 4'b1001 }: decoded = { 1'b0, 5'd04, 3'h1 };	// RD+
	{ 6'b101_001, 4'b1001 }: decoded = { 1'b0, 5'd05, 3'h1 };	// RD-/+
	// { 6'b101_001, 4'b1001 }: decoded = { 1'b0, 5'd05, 3'h1 };	// RD+
	{ 6'b011_001, 4'b1001 }: decoded = { 1'b0, 5'd06, 3'h1 };	// RD-/+
	// { 6'b011_001, 4'b1001 }: decoded = { 1'b0, 5'd06, 3'h1 };	// RD+
	{ 6'b111_000, 4'b1001 }: decoded = { 1'b0, 5'd07, 3'h1 };	// RD-
	{ 6'b000_111, 4'b1001 }: decoded = { 1'b0, 5'd07, 3'h1 };	// RD+
	//
	{ 6'b111_001, 4'b1001 }: decoded = { 1'b0, 5'd08, 3'h1 };	// RD-
	{ 6'b000_110, 4'b1001 }: decoded = { 1'b0, 5'd08, 3'h1 };	// RD+
	{ 6'b100_101, 4'b1001 }: decoded = { 1'b0, 5'd09, 3'h1 };	// RD-/+
	// { 6'b100_101, 4'b1001 }: decoded = { 1'b0, 5'd09, 3'h1 };	// RD+
	{ 6'b010_101, 4'b1001 }: decoded = { 1'b0, 5'd10, 3'h1 };	// RD-/+
	// { 6'b010_101, 4'b1001 }: decoded = { 1'b0, 5'd10, 3'h1 };	// RD+
	{ 6'b110_100, 4'b1001 }: decoded = { 1'b0, 5'd11, 3'h1 };	// RD-/+
	// { 6'b110_100, 4'b1001 }: decoded = { 1'b0, 5'd11, 3'h1 };	// RD+
	{ 6'b001_101, 4'b1001 }: decoded = { 1'b0, 5'd12, 3'h1 };	// RD-/+
	// { 6'b001_101, 4'b1001 }: decoded = { 1'b0, 5'd12, 3'h1 };	// RD+
	{ 6'b101_100, 4'b1001 }: decoded = { 1'b0, 5'd13, 3'h1 };	// RD-/+
	// { 6'b101_100, 4'b1001 }: decoded = { 1'b0, 5'd13, 3'h1 };	// RD+
	{ 6'b011_100, 4'b1001 }: decoded = { 1'b0, 5'd14, 3'h1 };	// RD-/+
	// { 6'b011_100, 4'b1001 }: decoded = { 1'b0, 5'd14, 3'h1 };	// RD+
	{ 6'b010_111, 4'b1001 }: decoded = { 1'b0, 5'd15, 3'h1 };	// RD-
	{ 6'b101_000, 4'b1001 }: decoded = { 1'b0, 5'd15, 3'h1 };	// RD+
	//
	{ 6'b011_011, 4'b1001 }: decoded = { 1'b0, 5'd16, 3'h1 };	// RD-
	{ 6'b100_100, 4'b1001 }: decoded = { 1'b0, 5'd16, 3'h1 };	// RD+
	{ 6'b100_011, 4'b1001 }: decoded = { 1'b0, 5'd17, 3'h1 };	// RD-
	// { 6'b100_011, 4'b1001 }: decoded = { 1'b0, 5'd17, 3'h1 };	// RD+
	{ 6'b010_011, 4'b1001 }: decoded = { 1'b0, 5'd18, 3'h1 };	// RD-
	// { 6'b010_011, 4'b1001 }: decoded = { 1'b0, 5'd18, 3'h1 };	// RD+
	{ 6'b110_010, 4'b1001 }: decoded = { 1'b0, 5'd19, 3'h1 };	// RD-
	// { 6'b110_010, 4'b1001 }: decoded = { 1'b0, 5'd19, 3'h1 };	// RD+
	{ 6'b001_011, 4'b1001 }: decoded = { 1'b0, 5'd20, 3'h1 };	// RD-
	// { 6'b001_011, 4'b1001 }: decoded = { 1'b0, 5'd20, 3'h1 };	// RD+
	{ 6'b101_010, 4'b1001 }: decoded = { 1'b0, 5'd21, 3'h1 };	// RD-
	// { 6'b101_010, 4'b1001 }: decoded = { 1'b0, 5'd21, 3'h1 };	// RD+
	{ 6'b011_010, 4'b1001 }: decoded = { 1'b0, 5'd22, 3'h1 };	// RD-
	// { 6'b011_010, 4'b1001 }: decoded = { 1'b0, 5'd22, 3'h1 };	// RD+
	{ 6'b111_010, 4'b1001 }: decoded = { 1'b0, 5'd23, 3'h1 };	// RD-
	{ 6'b000_101, 4'b1001 }: decoded = { 1'b0, 5'd23, 3'h1 };	// RD+
	//
	{ 6'b110_011, 4'b1001 }: decoded = { 1'b0, 5'd24, 3'h1 };	// RD-
	{ 6'b001_100, 4'b1001 }: decoded = { 1'b0, 5'd24, 3'h1 };	// RD+
	{ 6'b100_110, 4'b1001 }: decoded = { 1'b0, 5'd25, 3'h1 };	// RD-
	// { 6'b100_110, 4'b1001 }: decoded = { 1'b0, 5'd25, 3'h1 };	// RD+
	{ 6'b010_110, 4'b1001 }: decoded = { 1'b0, 5'd26, 3'h1 };	// RD-
	// { 6'b010_110, 4'b1001 }: decoded = { 1'b0, 5'd26, 3'h1 };	// RD+
	{ 6'b110_110, 4'b1001 }: decoded = { 1'b0, 5'd27, 3'h1 };	// RD-
	{ 6'b001_001, 4'b1001 }: decoded = { 1'b0, 5'd27, 3'h1 };	// RD+
	{ 6'b001_110, 4'b1001 }: decoded = { 1'b0, 5'd28, 3'h1 };	// RD-
	// { 6'b001_110, 4'b1001 }: decoded = { 1'b0, 5'd28, 3'h1 };	// RD+
	{ 6'b101_110, 4'b1001 }: decoded = { 1'b0, 5'd29, 3'h1 };	// RD-
	{ 6'b010_001, 4'b1001 }: decoded = { 1'b0, 5'd29, 3'h1 };	// RD+
	{ 6'b011_110, 4'b1001 }: decoded = { 1'b0, 5'd30, 3'h1 };	// RD-
	{ 6'b100_001, 4'b1001 }: decoded = { 1'b0, 5'd30, 3'h1 };	// RD+
	{ 6'b101_011, 4'b1001 }: decoded = { 1'b0, 5'd31, 3'h1 };	// RD-
	{ 6'b010_100, 4'b1001 }: decoded = { 1'b0, 5'd31, 3'h1 };	// RD+
	//
	//
	//
	{ 6'b100_111, 4'b0101 }: decoded = { 1'b0, 5'd00, 3'h2 };	// RD-
	{ 6'b011_000, 4'b0101 }: decoded = { 1'b0, 5'd00, 3'h2 };	// RD+
	{ 6'b011_101, 4'b0101 }: decoded = { 1'b0, 5'd01, 3'h2 };	// RD-
	{ 6'b100_010, 4'b0101 }: decoded = { 1'b0, 5'd01, 3'h2 };	// RD+
	{ 6'b101_101, 4'b0101 }: decoded = { 1'b0, 5'd02, 3'h2 };	// RD-
	{ 6'b010_010, 4'b0101 }: decoded = { 1'b0, 5'd02, 3'h2 };	// RD+
	{ 6'b110_001, 4'b0101 }: decoded = { 1'b0, 5'd03, 3'h2 };	// RD-
	// { 6'b110_001, 4'b0101 }: decoded = { 1'b0, 5'd03, 3'h2 };	// RD+
	{ 6'b110_101, 4'b0101 }: decoded = { 1'b0, 5'd04, 3'h2 };	// RD-
	{ 6'b001_010, 4'b0101 }: decoded = { 1'b0, 5'd04, 3'h2 };	// RD+
	{ 6'b101_001, 4'b0101 }: decoded = { 1'b0, 5'd05, 3'h2 };	// RD-
	// { 6'b101_001, 4'b0101 }: decoded = { 1'b0, 5'd05, 3'h2 };	// RD+
	{ 6'b011_001, 4'b0101 }: decoded = { 1'b0, 5'd06, 3'h2 };	// RD-
	// { 6'b011_001, 4'b0101 }: decoded = { 1'b0, 5'd06, 3'h2 };	// RD+
	{ 6'b111_000, 4'b0101 }: decoded = { 1'b0, 5'd07, 3'h2 };	// RD-
	{ 6'b000_111, 4'b0101 }: decoded = { 1'b0, 5'd07, 3'h2 };	// RD+
	//
	{ 6'b111_001, 4'b0101 }: decoded = { 1'b0, 5'd08, 3'h2 };	// RD-
	{ 6'b000_110, 4'b0101 }: decoded = { 1'b0, 5'd08, 3'h2 };	// RD+
	{ 6'b100_101, 4'b0101 }: decoded = { 1'b0, 5'd09, 3'h2 };	// RD-
	// { 6'b100_101, 4'b0101 }: decoded = { 1'b0, 5'd09, 3'h2 };	// RD+
	{ 6'b010_101, 4'b0101 }: decoded = { 1'b0, 5'd10, 3'h2 };	// RD-
	// { 6'b010_101, 4'b0101 }: decoded = { 1'b0, 5'd10, 3'h2 };	// RD+
	{ 6'b110_100, 4'b0101 }: decoded = { 1'b0, 5'd11, 3'h2 };	// RD-
	// { 6'b110_100, 4'b0101 }: decoded = { 1'b0, 5'd11, 3'h2 };	// RD+
	{ 6'b001_101, 4'b0101 }: decoded = { 1'b0, 5'd12, 3'h2 };	// RD-
	// { 6'b001_101, 4'b0101 }: decoded = { 1'b0, 5'd12, 3'h2 };	// RD+
	{ 6'b101_100, 4'b0101 }: decoded = { 1'b0, 5'd13, 3'h2 };	// RD-
	// { 6'b101_100, 4'b0101 }: decoded = { 1'b0, 5'd13, 3'h2 };	// RD+
	{ 6'b011_100, 4'b0101 }: decoded = { 1'b0, 5'd14, 3'h2 };	// RD-
	// { 6'b011_100, 4'b0101 }: decoded = { 1'b0, 5'd14, 3'h2 };	// RD+
	{ 6'b010_111, 4'b0101 }: decoded = { 1'b0, 5'd15, 3'h2 };	// RD-
	{ 6'b101_000, 4'b0101 }: decoded = { 1'b0, 5'd15, 3'h2 };	// RD+
	//
	{ 6'b011_011, 4'b0101 }: decoded = { 1'b0, 5'd16, 3'h2 };	// RD-
	{ 6'b100_100, 4'b0101 }: decoded = { 1'b0, 5'd16, 3'h2 };	// RD+
	{ 6'b100_011, 4'b0101 }: decoded = { 1'b0, 5'd17, 3'h2 };	// RD-
	// { 6'b100_011, 4'b0101 }: decoded = { 1'b0, 5'd17, 3'h2 };	// RD+
	{ 6'b010_011, 4'b0101 }: decoded = { 1'b0, 5'd18, 3'h2 };	// RD-
	// { 6'b010_011, 4'b0101 }: decoded = { 1'b0, 5'd18, 3'h2 };	// RD+
	{ 6'b110_010, 4'b0101 }: decoded = { 1'b0, 5'd19, 3'h2 };	// RD-
	// { 6'b110_010, 4'b0101 }: decoded = { 1'b0, 5'd19, 3'h2 };	// RD+
	{ 6'b001_011, 4'b0101 }: decoded = { 1'b0, 5'd20, 3'h2 };	// RD-
	// { 6'b001_011, 4'b0101 }: decoded = { 1'b0, 5'd20, 3'h2 };	// RD+
	{ 6'b101_010, 4'b0101 }: decoded = { 1'b0, 5'd21, 3'h2 };	// RD-
	// { 6'b101_010, 4'b0101 }: decoded = { 1'b0, 5'd21, 3'h2 };	// RD+
	{ 6'b011_010, 4'b0101 }: decoded = { 1'b0, 5'd22, 3'h2 };	// RD-
	// { 6'b011_010, 4'b0101 }: decoded = { 1'b0, 5'd22, 3'h2 };	// RD+
	{ 6'b111_010, 4'b0101 }: decoded = { 1'b0, 5'd23, 3'h2 };	// RD-
	{ 6'b000_101, 4'b0101 }: decoded = { 1'b0, 5'd23, 3'h2 };	// RD+
	//
	{ 6'b110_011, 4'b0101 }: decoded = { 1'b0, 5'd24, 3'h2 };	// RD-
	{ 6'b001_100, 4'b0101 }: decoded = { 1'b0, 5'd24, 3'h2 };	// RD+
	{ 6'b100_110, 4'b0101 }: decoded = { 1'b0, 5'd25, 3'h2 };	// RD-
	// { 6'b100_110, 4'b0101 }: decoded = { 1'b0, 5'd25, 3'h2 };	// RD+
	{ 6'b010_110, 4'b0101 }: decoded = { 1'b0, 5'd26, 3'h2 };	// RD-
	// { 6'b010_110, 4'b0101 }: decoded = { 1'b0, 5'd26, 3'h2 };	// RD+
	{ 6'b110_110, 4'b0101 }: decoded = { 1'b0, 5'd27, 3'h2 };	// RD-
	{ 6'b001_001, 4'b0101 }: decoded = { 1'b0, 5'd27, 3'h2 };	// RD+
	{ 6'b001_110, 4'b0101 }: decoded = { 1'b0, 5'd28, 3'h2 };	// RD-
	// { 6'b001_110, 4'b0101 }: decoded = { 1'b0, 5'd28, 3'h2 };	// RD+
	{ 6'b101_110, 4'b0101 }: decoded = { 1'b0, 5'd29, 3'h2 };	// RD-
	{ 6'b010_001, 4'b0101 }: decoded = { 1'b0, 5'd29, 3'h2 };	// RD+
	{ 6'b011_110, 4'b0101 }: decoded = { 1'b0, 5'd30, 3'h2 };	// RD-
	{ 6'b100_001, 4'b0101 }: decoded = { 1'b0, 5'd30, 3'h2 };	// RD+
	{ 6'b101_011, 4'b0101 }: decoded = { 1'b0, 5'd31, 3'h2 };	// RD-
	{ 6'b010_100, 4'b0101 }: decoded = { 1'b0, 5'd31, 3'h2 };	// RD+
	//
	//
	//
	{ 6'b100_111, 4'b0011 }: decoded = { 1'b0, 5'd00, 3'h3 };	// RD-
	{ 6'b011_000, 4'b1100 }: decoded = { 1'b0, 5'd00, 3'h3 };	// RD+
	{ 6'b011_101, 4'b0011 }: decoded = { 1'b0, 5'd01, 3'h3 };	// RD-
	{ 6'b100_010, 4'b1100 }: decoded = { 1'b0, 5'd01, 3'h3 };	// RD+
	{ 6'b101_101, 4'b0011 }: decoded = { 1'b0, 5'd02, 3'h3 };	// RD-
	{ 6'b010_010, 4'b1100 }: decoded = { 1'b0, 5'd02, 3'h3 };	// RD+
	{ 6'b110_001, 4'b1100 }: decoded = { 1'b0, 5'd03, 3'h3 };	// RD-
	{ 6'b110_001, 4'b0011 }: decoded = { 1'b0, 5'd03, 3'h3 };	// RD+
	{ 6'b110_101, 4'b0011 }: decoded = { 1'b0, 5'd04, 3'h3 };	// RD-
	{ 6'b001_010, 4'b1100 }: decoded = { 1'b0, 5'd04, 3'h3 };	// RD+
	{ 6'b101_001, 4'b1100 }: decoded = { 1'b0, 5'd05, 3'h3 };	// RD-
	{ 6'b101_001, 4'b0011 }: decoded = { 1'b0, 5'd05, 3'h3 };	// RD+
	{ 6'b011_001, 4'b1100 }: decoded = { 1'b0, 5'd06, 3'h3 };	// RD-
	{ 6'b011_001, 4'b0011 }: decoded = { 1'b0, 5'd06, 3'h3 };	// RD+
	{ 6'b111_000, 4'b1100 }: decoded = { 1'b0, 5'd07, 3'h3 };	// RD-
	{ 6'b000_111, 4'b0011 }: decoded = { 1'b0, 5'd07, 3'h3 };	// RD+
	//
	{ 6'b111_001, 4'b0011 }: decoded = { 1'b0, 5'd08, 3'h3 };	// RD-
	{ 6'b000_110, 4'b1100 }: decoded = { 1'b0, 5'd08, 3'h3 };	// RD+
	{ 6'b100_101, 4'b1100 }: decoded = { 1'b0, 5'd09, 3'h3 };	// RD-
	{ 6'b100_101, 4'b0011 }: decoded = { 1'b0, 5'd09, 3'h3 };	// RD+
	{ 6'b010_101, 4'b1100 }: decoded = { 1'b0, 5'd10, 3'h3 };	// RD-
	{ 6'b010_101, 4'b0011 }: decoded = { 1'b0, 5'd10, 3'h3 };	// RD+
	{ 6'b110_100, 4'b1100 }: decoded = { 1'b0, 5'd11, 3'h3 };	// RD-
	{ 6'b110_100, 4'b0011 }: decoded = { 1'b0, 5'd11, 3'h3 };	// RD+
	{ 6'b001_101, 4'b1100 }: decoded = { 1'b0, 5'd12, 3'h3 };	// RD-
	{ 6'b001_101, 4'b0011 }: decoded = { 1'b0, 5'd12, 3'h3 };	// RD+
	{ 6'b101_100, 4'b1100 }: decoded = { 1'b0, 5'd13, 3'h3 };	// RD-
	{ 6'b101_100, 4'b0011 }: decoded = { 1'b0, 5'd13, 3'h3 };	// RD+
	{ 6'b011_100, 4'b1100 }: decoded = { 1'b0, 5'd14, 3'h3 };	// RD-
	{ 6'b011_100, 4'b0011 }: decoded = { 1'b0, 5'd14, 3'h3 };	// RD+
	{ 6'b010_111, 4'b0011 }: decoded = { 1'b0, 5'd15, 3'h3 };	// RD-
	{ 6'b101_000, 4'b1100 }: decoded = { 1'b0, 5'd15, 3'h3 };	// RD+
	//
	{ 6'b011_011, 4'b0011 }: decoded = { 1'b0, 5'd16, 3'h3 };	// RD-
	{ 6'b100_100, 4'b1100 }: decoded = { 1'b0, 5'd16, 3'h3 };	// RD+
	{ 6'b100_011, 4'b1100 }: decoded = { 1'b0, 5'd17, 3'h3 };	// RD-
	{ 6'b100_011, 4'b0011 }: decoded = { 1'b0, 5'd17, 3'h3 };	// RD+
	{ 6'b010_011, 4'b1100 }: decoded = { 1'b0, 5'd18, 3'h3 };	// RD-
	{ 6'b010_011, 4'b0011 }: decoded = { 1'b0, 5'd18, 3'h3 };	// RD+
	{ 6'b110_010, 4'b1100 }: decoded = { 1'b0, 5'd19, 3'h3 };	// RD-
	{ 6'b110_010, 4'b0011 }: decoded = { 1'b0, 5'd19, 3'h3 };	// RD+
	{ 6'b001_011, 4'b1100 }: decoded = { 1'b0, 5'd20, 3'h3 };	// RD-
	{ 6'b001_011, 4'b0011 }: decoded = { 1'b0, 5'd20, 3'h3 };	// RD+
	{ 6'b101_010, 4'b1100 }: decoded = { 1'b0, 5'd21, 3'h3 };	// RD-
	{ 6'b101_010, 4'b0011 }: decoded = { 1'b0, 5'd21, 3'h3 };	// RD+
	{ 6'b011_010, 4'b1100 }: decoded = { 1'b0, 5'd22, 3'h3 };	// RD-
	{ 6'b011_010, 4'b0011 }: decoded = { 1'b0, 5'd22, 3'h3 };	// RD+
	{ 6'b111_010, 4'b0011 }: decoded = { 1'b0, 5'd23, 3'h3 };	// RD-
	{ 6'b000_101, 4'b1100 }: decoded = { 1'b0, 5'd23, 3'h3 };	// RD+
	//
	{ 6'b110_011, 4'b0011 }: decoded = { 1'b0, 5'd24, 3'h3 };	// RD-
	{ 6'b001_100, 4'b1100 }: decoded = { 1'b0, 5'd24, 3'h3 };	// RD+
	{ 6'b100_110, 4'b1100 }: decoded = { 1'b0, 5'd25, 3'h3 };	// RD-
	{ 6'b100_110, 4'b0011 }: decoded = { 1'b0, 5'd25, 3'h3 };	// RD+
	{ 6'b010_110, 4'b1100 }: decoded = { 1'b0, 5'd26, 3'h3 };	// RD-
	{ 6'b010_110, 4'b0011 }: decoded = { 1'b0, 5'd26, 3'h3 };	// RD+
	{ 6'b110_110, 4'b0011 }: decoded = { 1'b0, 5'd27, 3'h3 };	// RD-
	{ 6'b001_001, 4'b1100 }: decoded = { 1'b0, 5'd27, 3'h3 };	// RD+
	{ 6'b001_110, 4'b1100 }: decoded = { 1'b0, 5'd28, 3'h3 };	// RD-
	{ 6'b001_110, 4'b0011 }: decoded = { 1'b0, 5'd28, 3'h3 };	// RD+
	{ 6'b101_110, 4'b0011 }: decoded = { 1'b0, 5'd29, 3'h3 };	// RD-
	{ 6'b010_001, 4'b1100 }: decoded = { 1'b0, 5'd29, 3'h3 };	// RD+
	{ 6'b011_110, 4'b0011 }: decoded = { 1'b0, 5'd30, 3'h3 };	// RD-
	{ 6'b100_001, 4'b1100 }: decoded = { 1'b0, 5'd30, 3'h3 };	// RD+
	{ 6'b101_011, 4'b0011 }: decoded = { 1'b0, 5'd31, 3'h3 };	// RD-
	{ 6'b010_100, 4'b1100 }: decoded = { 1'b0, 5'd31, 3'h3 };	// RD+
	//
	//
	//
	{ 6'b100_111, 4'b0010 }: decoded = { 1'b0, 5'd00, 3'h4 };	// RD-
	{ 6'b011_000, 4'b1101 }: decoded = { 1'b0, 5'd00, 3'h4 };	// RD+
	{ 6'b011_101, 4'b0010 }: decoded = { 1'b0, 5'd01, 3'h4 };	// RD-
	{ 6'b100_010, 4'b1101 }: decoded = { 1'b0, 5'd01, 3'h4 };	// RD+
	{ 6'b101_101, 4'b0010 }: decoded = { 1'b0, 5'd02, 3'h4 };	// RD-
	{ 6'b010_010, 4'b1101 }: decoded = { 1'b0, 5'd02, 3'h4 };	// RD+
	{ 6'b110_001, 4'b1101 }: decoded = { 1'b0, 5'd03, 3'h4 };	// RD-
	{ 6'b110_001, 4'b0010 }: decoded = { 1'b0, 5'd03, 3'h4 };	// RD+
	{ 6'b110_101, 4'b0010 }: decoded = { 1'b0, 5'd04, 3'h4 };	// RD-
	{ 6'b001_010, 4'b1101 }: decoded = { 1'b0, 5'd04, 3'h4 };	// RD+
	{ 6'b101_001, 4'b1101 }: decoded = { 1'b0, 5'd05, 3'h4 };	// RD-
	{ 6'b101_001, 4'b0010 }: decoded = { 1'b0, 5'd05, 3'h4 };	// RD+
	{ 6'b011_001, 4'b1101 }: decoded = { 1'b0, 5'd06, 3'h4 };	// RD-
	{ 6'b011_001, 4'b0010 }: decoded = { 1'b0, 5'd06, 3'h4 };	// RD+
	{ 6'b111_000, 4'b1101 }: decoded = { 1'b0, 5'd07, 3'h4 };	// RD-
	{ 6'b000_111, 4'b0010 }: decoded = { 1'b0, 5'd07, 3'h4 };	// RD+
	//
	{ 6'b111_001, 4'b0010 }: decoded = { 1'b0, 5'd08, 3'h4 };	// RD-
	{ 6'b000_110, 4'b1101 }: decoded = { 1'b0, 5'd08, 3'h4 };	// RD+
	{ 6'b100_101, 4'b1101 }: decoded = { 1'b0, 5'd09, 3'h4 };	// RD-
	{ 6'b100_101, 4'b0010 }: decoded = { 1'b0, 5'd09, 3'h4 };	// RD+
	{ 6'b010_101, 4'b1101 }: decoded = { 1'b0, 5'd10, 3'h4 };	// RD-
	{ 6'b010_101, 4'b0010 }: decoded = { 1'b0, 5'd10, 3'h4 };	// RD+
	{ 6'b110_100, 4'b1101 }: decoded = { 1'b0, 5'd11, 3'h4 };	// RD-
	{ 6'b110_100, 4'b0010 }: decoded = { 1'b0, 5'd11, 3'h4 };	// RD+
	{ 6'b001_101, 4'b1101 }: decoded = { 1'b0, 5'd12, 3'h4 };	// RD-
	{ 6'b001_101, 4'b0010 }: decoded = { 1'b0, 5'd12, 3'h4 };	// RD+
	{ 6'b101_100, 4'b1101 }: decoded = { 1'b0, 5'd13, 3'h4 };	// RD-
	{ 6'b101_100, 4'b0010 }: decoded = { 1'b0, 5'd13, 3'h4 };	// RD+
	{ 6'b011_100, 4'b1101 }: decoded = { 1'b0, 5'd14, 3'h4 };	// RD-
	{ 6'b011_100, 4'b0010 }: decoded = { 1'b0, 5'd14, 3'h4 };	// RD+
	{ 6'b010_111, 4'b0010 }: decoded = { 1'b0, 5'd15, 3'h4 };	// RD-
	{ 6'b101_000, 4'b1101 }: decoded = { 1'b0, 5'd15, 3'h4 };	// RD+
	//
	{ 6'b011_011, 4'b0010 }: decoded = { 1'b0, 5'd16, 3'h4 };	// RD-
	{ 6'b100_100, 4'b1101 }: decoded = { 1'b0, 5'd16, 3'h4 };	// RD+
	{ 6'b100_011, 4'b1101 }: decoded = { 1'b0, 5'd17, 3'h4 };	// RD-
	{ 6'b100_011, 4'b0010 }: decoded = { 1'b0, 5'd17, 3'h4 };	// RD+
	{ 6'b010_011, 4'b1101 }: decoded = { 1'b0, 5'd18, 3'h4 };	// RD-
	{ 6'b010_011, 4'b0010 }: decoded = { 1'b0, 5'd18, 3'h4 };	// RD+
	{ 6'b110_010, 4'b1101 }: decoded = { 1'b0, 5'd19, 3'h4 };	// RD-
	{ 6'b110_010, 4'b0010 }: decoded = { 1'b0, 5'd19, 3'h4 };	// RD+
	{ 6'b001_011, 4'b1101 }: decoded = { 1'b0, 5'd20, 3'h4 };	// RD-
	{ 6'b001_011, 4'b0010 }: decoded = { 1'b0, 5'd20, 3'h4 };	// RD+
	{ 6'b101_010, 4'b1101 }: decoded = { 1'b0, 5'd21, 3'h4 };	// RD-
	{ 6'b101_010, 4'b0010 }: decoded = { 1'b0, 5'd21, 3'h4 };	// RD+
	{ 6'b011_010, 4'b1101 }: decoded = { 1'b0, 5'd22, 3'h4 };	// RD-
	{ 6'b011_010, 4'b0010 }: decoded = { 1'b0, 5'd22, 3'h4 };	// RD+
	{ 6'b111_010, 4'b0010 }: decoded = { 1'b0, 5'd23, 3'h4 };	// RD-
	{ 6'b000_101, 4'b1101 }: decoded = { 1'b0, 5'd23, 3'h4 };	// RD+
	//
	{ 6'b110_011, 4'b0010 }: decoded = { 1'b0, 5'd24, 3'h4 };	// RD-
	{ 6'b001_100, 4'b1101 }: decoded = { 1'b0, 5'd24, 3'h4 };	// RD+
	{ 6'b100_110, 4'b1101 }: decoded = { 1'b0, 5'd25, 3'h4 };	// RD-
	{ 6'b100_110, 4'b0010 }: decoded = { 1'b0, 5'd25, 3'h4 };	// RD+
	{ 6'b010_110, 4'b1101 }: decoded = { 1'b0, 5'd26, 3'h4 };	// RD-
	{ 6'b010_110, 4'b0010 }: decoded = { 1'b0, 5'd26, 3'h4 };	// RD+
	{ 6'b110_110, 4'b0010 }: decoded = { 1'b0, 5'd27, 3'h4 };	// RD-
	{ 6'b001_001, 4'b1101 }: decoded = { 1'b0, 5'd27, 3'h4 };	// RD+
	{ 6'b001_110, 4'b1101 }: decoded = { 1'b0, 5'd28, 3'h4 };	// RD-
	{ 6'b001_110, 4'b0010 }: decoded = { 1'b0, 5'd28, 3'h4 };	// RD+
	{ 6'b101_110, 4'b0010 }: decoded = { 1'b0, 5'd29, 3'h4 };	// RD-
	{ 6'b010_001, 4'b1101 }: decoded = { 1'b0, 5'd29, 3'h4 };	// RD+
	{ 6'b011_110, 4'b0010 }: decoded = { 1'b0, 5'd30, 3'h4 };	// RD-
	{ 6'b100_001, 4'b1101 }: decoded = { 1'b0, 5'd30, 3'h4 };	// RD+
	{ 6'b101_011, 4'b0010 }: decoded = { 1'b0, 5'd31, 3'h4 };	// RD-
	{ 6'b010_100, 4'b1101 }: decoded = { 1'b0, 5'd31, 3'h4 };	// RD+
	//
	//
	//
	{ 6'b100_111, 4'b1010 }: decoded = { 1'b0, 5'd00, 3'h5 };	// RD-
	{ 6'b011_000, 4'b1010 }: decoded = { 1'b0, 5'd00, 3'h5 };	// RD+
	{ 6'b011_101, 4'b1010 }: decoded = { 1'b0, 5'd01, 3'h5 };	// RD-
	{ 6'b100_010, 4'b1010 }: decoded = { 1'b0, 5'd01, 3'h5 };	// RD+
	{ 6'b101_101, 4'b1010 }: decoded = { 1'b0, 5'd02, 3'h5 };	// RD-
	{ 6'b010_010, 4'b1010 }: decoded = { 1'b0, 5'd02, 3'h5 };	// RD+
	{ 6'b110_001, 4'b1010 }: decoded = { 1'b0, 5'd03, 3'h5 };	// RD-
	// { 6'b110_001, 4'b1010 }: decoded = { 1'b0, 5'd03, 3'h5 };	// RD+
	{ 6'b110_101, 4'b1010 }: decoded = { 1'b0, 5'd04, 3'h5 };	// RD-
	{ 6'b001_010, 4'b1010 }: decoded = { 1'b0, 5'd04, 3'h5 };	// RD+
	{ 6'b101_001, 4'b1010 }: decoded = { 1'b0, 5'd05, 3'h5 };	// RD-
	// { 6'b101_001, 4'b1010 }: decoded = { 1'b0, 5'd05, 3'h5 };	// RD+
	{ 6'b011_001, 4'b1010 }: decoded = { 1'b0, 5'd06, 3'h5 };	// RD-
	// { 6'b011_001, 4'b1010 }: decoded = { 1'b0, 5'd06, 3'h5 };	// RD+
	{ 6'b111_000, 4'b1010 }: decoded = { 1'b0, 5'd07, 3'h5 };	// RD-
	{ 6'b000_111, 4'b1010 }: decoded = { 1'b0, 5'd07, 3'h5 };	// RD+
	//
	{ 6'b111_001, 4'b1010 }: decoded = { 1'b0, 5'd08, 3'h5 };	// RD-
	{ 6'b000_110, 4'b1010 }: decoded = { 1'b0, 5'd08, 3'h5 };	// RD+
	{ 6'b100_101, 4'b1010 }: decoded = { 1'b0, 5'd09, 3'h5 };	// RD-
	// { 6'b100_101, 4'b1010 }: decoded = { 1'b0, 5'd09, 3'h5 };	// RD+
	{ 6'b010_101, 4'b1010 }: decoded = { 1'b0, 5'd10, 3'h5 };	// RD-
	// { 6'b010_101, 4'b1010 }: decoded = { 1'b0, 5'd10, 3'h5 };	// RD+
	{ 6'b110_100, 4'b1010 }: decoded = { 1'b0, 5'd11, 3'h5 };	// RD-
	// { 6'b110_100, 4'b1010 }: decoded = { 1'b0, 5'd11, 3'h5 };	// RD+
	{ 6'b001_101, 4'b1010 }: decoded = { 1'b0, 5'd12, 3'h5 };	// RD-
	// { 6'b001_101, 4'b1010 }: decoded = { 1'b0, 5'd12, 3'h5 };	// RD+
	{ 6'b101_100, 4'b1010 }: decoded = { 1'b0, 5'd13, 3'h5 };	// RD-
	// { 6'b101_100, 4'b1010 }: decoded = { 1'b0, 5'd13, 3'h5 };	// RD+
	{ 6'b011_100, 4'b1010 }: decoded = { 1'b0, 5'd14, 3'h5 };	// RD-
	// { 6'b011_100, 4'b1010 }: decoded = { 1'b0, 5'd14, 3'h5 };	// RD+
	{ 6'b010_111, 4'b1010 }: decoded = { 1'b0, 5'd15, 3'h5 };	// RD-
	{ 6'b101_000, 4'b1010 }: decoded = { 1'b0, 5'd15, 3'h5 };	// RD+
	//
	{ 6'b011_011, 4'b1010 }: decoded = { 1'b0, 5'd16, 3'h5 };	// RD-
	{ 6'b100_100, 4'b1010 }: decoded = { 1'b0, 5'd16, 3'h5 };	// RD+
	{ 6'b100_011, 4'b1010 }: decoded = { 1'b0, 5'd17, 3'h5 };	// RD-
	// { 6'b100_011, 4'b1010 }: decoded = { 1'b0, 5'd17, 3'h5 };	// RD+
	{ 6'b010_011, 4'b1010 }: decoded = { 1'b0, 5'd18, 3'h5 };	// RD-
	// { 6'b010_011, 4'b1010 }: decoded = { 1'b0, 5'd18, 3'h5 };	// RD+
	{ 6'b110_010, 4'b1010 }: decoded = { 1'b0, 5'd19, 3'h5 };	// RD-
	// { 6'b110_010, 4'b1010 }: decoded = { 1'b0, 5'd19, 3'h5 };	// RD+
	{ 6'b001_011, 4'b1010 }: decoded = { 1'b0, 5'd20, 3'h5 };	// RD-
	// { 6'b001_011, 4'b1010 }: decoded = { 1'b0, 5'd20, 3'h5 };	// RD+
	{ 6'b101_010, 4'b1010 }: decoded = { 1'b0, 5'd21, 3'h5 };	// RD-
	// { 6'b101_010, 4'b1010 }: decoded = { 1'b0, 5'd21, 3'h5 };	// RD+
	{ 6'b011_010, 4'b1010 }: decoded = { 1'b0, 5'd22, 3'h5 };	// RD-
	// { 6'b011_010, 4'b1010 }: decoded = { 1'b0, 5'd22, 3'h5 };	// RD+
	{ 6'b111_010, 4'b1010 }: decoded = { 1'b0, 5'd23, 3'h5 };	// RD-
	{ 6'b000_101, 4'b1010 }: decoded = { 1'b0, 5'd23, 3'h5 };	// RD+
	//
	{ 6'b110_011, 4'b1010 }: decoded = { 1'b0, 5'd24, 3'h5 };	// RD-
	{ 6'b001_100, 4'b1010 }: decoded = { 1'b0, 5'd24, 3'h5 };	// RD+
	{ 6'b100_110, 4'b1010 }: decoded = { 1'b0, 5'd25, 3'h5 };	// RD-
	// { 6'b100_110, 4'b1010 }: decoded = { 1'b0, 5'd25, 3'h5 };	// RD+
	{ 6'b010_110, 4'b1010 }: decoded = { 1'b0, 5'd26, 3'h5 };	// RD-
	// { 6'b010_110, 4'b1010 }: decoded = { 1'b0, 5'd26, 3'h5 };	// RD+
	{ 6'b110_110, 4'b1010 }: decoded = { 1'b0, 5'd27, 3'h5 };	// RD-
	{ 6'b001_001, 4'b1010 }: decoded = { 1'b0, 5'd27, 3'h5 };	// RD+
	{ 6'b001_110, 4'b1010 }: decoded = { 1'b0, 5'd28, 3'h5 };	// RD-
	// { 6'b001_110, 4'b1010 }: decoded = { 1'b0, 5'd28, 3'h5 };	// RD+
	{ 6'b101_110, 4'b1010 }: decoded = { 1'b0, 5'd29, 3'h5 };	// RD-
	{ 6'b010_001, 4'b1010 }: decoded = { 1'b0, 5'd29, 3'h5 };	// RD+
	{ 6'b011_110, 4'b1010 }: decoded = { 1'b0, 5'd30, 3'h5 };	// RD-
	{ 6'b100_001, 4'b1010 }: decoded = { 1'b0, 5'd30, 3'h5 };	// RD+
	{ 6'b101_011, 4'b1010 }: decoded = { 1'b0, 5'd31, 3'h5 };	// RD-
	{ 6'b010_100, 4'b1010 }: decoded = { 1'b0, 5'd31, 3'h5 };	// RD+
	//
	//
	//
	{ 6'b100_111, 4'b0110 }: decoded = { 1'b0, 5'd00, 3'h6 };	// RD-
	{ 6'b011_000, 4'b0110 }: decoded = { 1'b0, 5'd00, 3'h6 };	// RD+
	{ 6'b011_101, 4'b0110 }: decoded = { 1'b0, 5'd01, 3'h6 };	// RD-
	{ 6'b100_010, 4'b0110 }: decoded = { 1'b0, 5'd01, 3'h6 };	// RD+
	{ 6'b101_101, 4'b0110 }: decoded = { 1'b0, 5'd02, 3'h6 };	// RD-
	{ 6'b010_010, 4'b0110 }: decoded = { 1'b0, 5'd02, 3'h6 };	// RD+
	{ 6'b110_001, 4'b0110 }: decoded = { 1'b0, 5'd03, 3'h6 };	// RD-
	// { 6'b110_001, 4'b0110 }: decoded = { 1'b0, 5'd03, 3'h6 };	// RD+
	{ 6'b110_101, 4'b0110 }: decoded = { 1'b0, 5'd04, 3'h6 };	// RD-
	{ 6'b001_010, 4'b0110 }: decoded = { 1'b0, 5'd04, 3'h6 };	// RD+
	{ 6'b101_001, 4'b0110 }: decoded = { 1'b0, 5'd05, 3'h6 };	// RD-
	// { 6'b101_001, 4'b0110 }: decoded = { 1'b0, 5'd05, 3'h6 };	// RD+
	{ 6'b011_001, 4'b0110 }: decoded = { 1'b0, 5'd06, 3'h6 };	// RD-
	// { 6'b011_001, 4'b0110 }: decoded = { 1'b0, 5'd06, 3'h6 };	// RD+
	{ 6'b111_000, 4'b0110 }: decoded = { 1'b0, 5'd07, 3'h6 };	// RD-
	{ 6'b000_111, 4'b0110 }: decoded = { 1'b0, 5'd07, 3'h6 };	// RD+
	//
	{ 6'b111_001, 4'b0110 }: decoded = { 1'b0, 5'd08, 3'h6 };	// RD-
	{ 6'b000_110, 4'b0110 }: decoded = { 1'b0, 5'd08, 3'h6 };	// RD+
	{ 6'b100_101, 4'b0110 }: decoded = { 1'b0, 5'd09, 3'h6 };	// RD-
	// { 6'b100_101, 4'b0110 }: decoded = { 1'b0, 5'd09, 3'h6 };	// RD+
	{ 6'b010_101, 4'b0110 }: decoded = { 1'b0, 5'd10, 3'h6 };	// RD-
	// { 6'b010_101, 4'b0110 }: decoded = { 1'b0, 5'd10, 3'h6 };	// RD+
	{ 6'b110_100, 4'b0110 }: decoded = { 1'b0, 5'd11, 3'h6 };	// RD-
	// { 6'b110_100, 4'b0110 }: decoded = { 1'b0, 5'd11, 3'h6 };	// RD+
	{ 6'b001_101, 4'b0110 }: decoded = { 1'b0, 5'd12, 3'h6 };	// RD-
	// { 6'b001_101, 4'b0110 }: decoded = { 1'b0, 5'd12, 3'h6 };	// RD+
	{ 6'b101_100, 4'b0110 }: decoded = { 1'b0, 5'd13, 3'h6 };	// RD-
	// { 6'b101_100, 4'b0110 }: decoded = { 1'b0, 5'd13, 3'h6 };	// RD+
	{ 6'b011_100, 4'b0110 }: decoded = { 1'b0, 5'd14, 3'h6 };	// RD-
	// { 6'b011_100, 4'b0110 }: decoded = { 1'b0, 5'd14, 3'h6 };	// RD+
	{ 6'b010_111, 4'b0110 }: decoded = { 1'b0, 5'd15, 3'h6 };	// RD-
	{ 6'b101_000, 4'b0110 }: decoded = { 1'b0, 5'd15, 3'h6 };	// RD+
	//
	{ 6'b011_011, 4'b0110 }: decoded = { 1'b0, 5'd16, 3'h6 };	// RD-
	{ 6'b100_100, 4'b0110 }: decoded = { 1'b0, 5'd16, 3'h6 };	// RD+
	{ 6'b100_011, 4'b0110 }: decoded = { 1'b0, 5'd17, 3'h6 };	// RD-
	// { 6'b100_011, 4'b0110 }: decoded = { 1'b0, 5'd17, 3'h6 };	// RD+
	{ 6'b010_011, 4'b0110 }: decoded = { 1'b0, 5'd18, 3'h6 };	// RD-
	// { 6'b010_011, 4'b0110 }: decoded = { 1'b0, 5'd18, 3'h6 };	// RD+
	{ 6'b110_010, 4'b0110 }: decoded = { 1'b0, 5'd19, 3'h6 };	// RD-
	// { 6'b110_010, 4'b0110 }: decoded = { 1'b0, 5'd19, 3'h6 };	// RD+
	{ 6'b001_011, 4'b0110 }: decoded = { 1'b0, 5'd20, 3'h6 };	// RD-
	// { 6'b001_011, 4'b0110 }: decoded = { 1'b0, 5'd20, 3'h6 };	// RD+
	{ 6'b101_010, 4'b0110 }: decoded = { 1'b0, 5'd21, 3'h6 };	// RD-
	// { 6'b101_010, 4'b0110 }: decoded = { 1'b0, 5'd21, 3'h6 };	// RD+
	{ 6'b011_010, 4'b0110 }: decoded = { 1'b0, 5'd22, 3'h6 };	// RD-
	// { 6'b011_010, 4'b0110 }: decoded = { 1'b0, 5'd22, 3'h6 };	// RD+
	{ 6'b111_010, 4'b0110 }: decoded = { 1'b0, 5'd23, 3'h6 };	// RD-
	{ 6'b000_101, 4'b0110 }: decoded = { 1'b0, 5'd23, 3'h6 };	// RD+
	//
	{ 6'b110_011, 4'b0110 }: decoded = { 1'b0, 5'd24, 3'h6 };	// RD-
	{ 6'b001_100, 4'b0110 }: decoded = { 1'b0, 5'd24, 3'h6 };	// RD+
	{ 6'b100_110, 4'b0110 }: decoded = { 1'b0, 5'd25, 3'h6 };	// RD-
	// { 6'b100_110, 4'b0110 }: decoded = { 1'b0, 5'd25, 3'h6 };	// RD+
	{ 6'b010_110, 4'b0110 }: decoded = { 1'b0, 5'd26, 3'h6 };	// RD-
	// { 6'b010_110, 4'b0110 }: decoded = { 1'b0, 5'd26, 3'h6 };	// RD+
	{ 6'b110_110, 4'b0110 }: decoded = { 1'b0, 5'd27, 3'h6 };	// RD-
	{ 6'b001_001, 4'b0110 }: decoded = { 1'b0, 5'd27, 3'h6 };	// RD+
	{ 6'b001_110, 4'b0110 }: decoded = { 1'b0, 5'd28, 3'h6 };	// RD-
	// { 6'b001_110, 4'b0110 }: decoded = { 1'b0, 5'd28, 3'h6 };	// RD+
	{ 6'b101_110, 4'b0110 }: decoded = { 1'b0, 5'd29, 3'h6 };	// RD-
	{ 6'b010_001, 4'b0110 }: decoded = { 1'b0, 5'd29, 3'h6 };	// RD+
	{ 6'b011_110, 4'b0110 }: decoded = { 1'b0, 5'd30, 3'h6 };	// RD-
	{ 6'b100_001, 4'b0110 }: decoded = { 1'b0, 5'd30, 3'h6 };	// RD+
	{ 6'b101_011, 4'b0110 }: decoded = { 1'b0, 5'd31, 3'h6 };	// RD-
	{ 6'b010_100, 4'b0110 }: decoded = { 1'b0, 5'd31, 3'h6 };	// RD+
	//
	//
	//
	{ 6'b100_111, 4'b0001 }: decoded = { 1'b0, 5'd00, 3'h7 };	// RD-
	{ 6'b011_000, 4'b1110 }: decoded = { 1'b0, 5'd00, 3'h7 };	// RD+
	{ 6'b011_101, 4'b0001 }: decoded = { 1'b0, 5'd01, 3'h7 };	// RD-
	{ 6'b100_010, 4'b1110 }: decoded = { 1'b0, 5'd01, 3'h7 };	// RD+
	{ 6'b101_101, 4'b0001 }: decoded = { 1'b0, 5'd02, 3'h7 };	// RD-
	{ 6'b010_010, 4'b1110 }: decoded = { 1'b0, 5'd02, 3'h7 };	// RD+
	{ 6'b110_001, 4'b1110 }: decoded = { 1'b0, 5'd03, 3'h7 };	// RD-
	{ 6'b110_001, 4'b0001 }: decoded = { 1'b0, 5'd03, 3'h7 };	// RD+
	{ 6'b110_101, 4'b0001 }: decoded = { 1'b0, 5'd04, 3'h7 };	// RD-
	{ 6'b001_010, 4'b1110 }: decoded = { 1'b0, 5'd04, 3'h7 };	// RD+
	{ 6'b101_001, 4'b1110 }: decoded = { 1'b0, 5'd05, 3'h7 };	// RD-
	{ 6'b101_001, 4'b0001 }: decoded = { 1'b0, 5'd05, 3'h7 };	// RD+
	{ 6'b011_001, 4'b1110 }: decoded = { 1'b0, 5'd06, 3'h7 };	// RD-
	{ 6'b011_001, 4'b0001 }: decoded = { 1'b0, 5'd06, 3'h7 };	// RD+
	{ 6'b111_000, 4'b1110 }: decoded = { 1'b0, 5'd07, 3'h7 };	// RD-
	{ 6'b000_111, 4'b0001 }: decoded = { 1'b0, 5'd07, 3'h7 };	// RD+
	//
	{ 6'b111_001, 4'b0001 }: decoded = { 1'b0, 5'd08, 3'h7 };	// RD-
	{ 6'b000_110, 4'b1110 }: decoded = { 1'b0, 5'd08, 3'h7 };	// RD+
	{ 6'b100_101, 4'b1110 }: decoded = { 1'b0, 5'd09, 3'h7 };	// RD-
	{ 6'b100_101, 4'b0001 }: decoded = { 1'b0, 5'd09, 3'h7 };	// RD+
	{ 6'b010_101, 4'b1110 }: decoded = { 1'b0, 5'd10, 3'h7 };	// RD-
	{ 6'b010_101, 4'b0001 }: decoded = { 1'b0, 5'd10, 3'h7 };	// RD+
	{ 6'b110_100, 4'b1110 }: decoded = { 1'b0, 5'd11, 3'h7 };	// RD-
	{ 6'b110_100, 4'b1000 }: decoded = { 1'b0, 5'd11, 3'h7 };	// RD+
	{ 6'b001_101, 4'b1110 }: decoded = { 1'b0, 5'd12, 3'h7 };	// RD-
	{ 6'b001_101, 4'b0001 }: decoded = { 1'b0, 5'd12, 3'h7 };	// RD+
	{ 6'b101_100, 4'b1110 }: decoded = { 1'b0, 5'd13, 3'h7 };	// RD-
	{ 6'b101_100, 4'b1000 }: decoded = { 1'b0, 5'd13, 3'h7 };	// RD+
	{ 6'b011_100, 4'b1110 }: decoded = { 1'b0, 5'd14, 3'h7 };	// RD-
	{ 6'b011_100, 4'b1000 }: decoded = { 1'b0, 5'd14, 3'h7 };	// RD+
	{ 6'b010_111, 4'b0001 }: decoded = { 1'b0, 5'd15, 3'h7 };	// RD-
	{ 6'b101_000, 4'b1110 }: decoded = { 1'b0, 5'd15, 3'h7 };	// RD+
	//
	{ 6'b011_011, 4'b0001 }: decoded = { 1'b0, 5'd16, 3'h7 };	// RD-
	{ 6'b100_100, 4'b1110 }: decoded = { 1'b0, 5'd16, 3'h7 };	// RD+
	{ 6'b100_011, 4'b0111 }: decoded = { 1'b0, 5'd17, 3'h7 };	// RD-
	{ 6'b100_011, 4'b0001 }: decoded = { 1'b0, 5'd17, 3'h7 };	// RD+
	{ 6'b010_011, 4'b0111 }: decoded = { 1'b0, 5'd18, 3'h7 };	// RD-
	{ 6'b010_011, 4'b0001 }: decoded = { 1'b0, 5'd18, 3'h7 };	// RD+
	{ 6'b110_010, 4'b1110 }: decoded = { 1'b0, 5'd19, 3'h7 };	// RD-
	{ 6'b110_010, 4'b0001 }: decoded = { 1'b0, 5'd19, 3'h7 };	// RD+
	{ 6'b001_011, 4'b0111 }: decoded = { 1'b0, 5'd20, 3'h7 };	// RD-
	{ 6'b001_011, 4'b0001 }: decoded = { 1'b0, 5'd20, 3'h7 };	// RD+
	{ 6'b101_010, 4'b1110 }: decoded = { 1'b0, 5'd21, 3'h7 };	// RD-
	{ 6'b101_010, 4'b0001 }: decoded = { 1'b0, 5'd21, 3'h7 };	// RD+
	{ 6'b011_010, 4'b1110 }: decoded = { 1'b0, 5'd22, 3'h7 };	// RD-
	{ 6'b011_010, 4'b0001 }: decoded = { 1'b0, 5'd22, 3'h7 };	// RD+
	{ 6'b111_010, 4'b0001 }: decoded = { 1'b0, 5'd23, 3'h7 };	// RD-
	{ 6'b000_101, 4'b1110 }: decoded = { 1'b0, 5'd23, 3'h7 };	// RD+
	//
	{ 6'b110_011, 4'b0001 }: decoded = { 1'b0, 5'd24, 3'h7 };	// RD-
	{ 6'b001_100, 4'b1110 }: decoded = { 1'b0, 5'd24, 3'h7 };	// RD+
	{ 6'b100_110, 4'b1110 }: decoded = { 1'b0, 5'd25, 3'h7 };	// RD-
	{ 6'b100_110, 4'b0001 }: decoded = { 1'b0, 5'd25, 3'h7 };	// RD+
	{ 6'b010_110, 4'b1110 }: decoded = { 1'b0, 5'd26, 3'h7 };	// RD-
	{ 6'b010_110, 4'b0001 }: decoded = { 1'b0, 5'd26, 3'h7 };	// RD+
	{ 6'b110_110, 4'b0001 }: decoded = { 1'b0, 5'd27, 3'h7 };	// RD-
	{ 6'b001_001, 4'b1110 }: decoded = { 1'b0, 5'd27, 3'h7 };	// RD+
	{ 6'b001_110, 4'b1110 }: decoded = { 1'b0, 5'd28, 3'h7 };	// RD-
	{ 6'b001_110, 4'b0001 }: decoded = { 1'b0, 5'd28, 3'h7 };	// RD+
	{ 6'b101_110, 4'b0001 }: decoded = { 1'b0, 5'd29, 3'h7 };	// RD-
	{ 6'b010_001, 4'b1110 }: decoded = { 1'b0, 5'd29, 3'h7 };	// RD+
	{ 6'b011_110, 4'b0001 }: decoded = { 1'b0, 5'd30, 3'h7 };	// RD-
	{ 6'b100_001, 4'b1110 }: decoded = { 1'b0, 5'd30, 3'h7 };	// RD+
	{ 6'b101_011, 4'b0001 }: decoded = { 1'b0, 5'd31, 3'h7 };	// RD-
	{ 6'b010_100, 4'b1110 }: decoded = { 1'b0, 5'd31, 3'h7 };	// RD+
	//
	{ 6'b001_111, 4'b0011 }: decoded = { 1'b1, 5'd28, 3'h3 };	// RD-
	{ 6'b110_000, 4'b1100 }: decoded = { 1'b1, 5'd28, 3'h3 };	// RD+
	{ 6'b001_111, 4'b1010 }: decoded = { 1'b1, 5'd28, 3'h5 };	// RD-
	{ 6'b110_000, 4'b0101 }: decoded = { 1'b1, 5'd28, 3'h5 };	// RD+
	//
	default: decoded = { 1'b1, 8'hff };
	endcase

	assign M_DATA = { decoded[8], decoded[2:0], decoded[7:3] };

////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////
//
// Formal properties
// {{{
////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////
`ifdef	FORMAL
	(* keep *) wire	[4:0]	Dx = decoded[8:3];
	(* keep *) wire	[2:0]	Dy = decoded[2:0];
`endif
// }}}
endmodule
